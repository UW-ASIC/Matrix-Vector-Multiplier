** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/TIAs/optimization_temp/TIA_optimization/TIA_temp_opt/tb/TIA_TO_test_tb.sch
**.subckt TIA_TO_test_tb
*  x1 -  TIA  IS MISSING !!!!
I0 net1 Iin 1m
V1 net2 GND 3
V2 net3 GND 3
**** begin user architecture code

.op


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
