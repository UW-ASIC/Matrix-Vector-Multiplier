** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/TIAs/OpAmp_temp_opt/tb/OpAmp_TO_slew_rate_tb.sch
**.subckt OpAmp_TO_slew_rate_tb
**.ends
.end
