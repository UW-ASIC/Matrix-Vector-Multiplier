** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/TIAs/TIA_LowNoise/tb/TIA_LN_power_consumption_tb.sch
**.subckt TIA_LN_power_consumption_tb
*  x1 -  TIA  IS MISSING !!!!
I0 net1 Iin DC 1u
V1 net2 GND DC 3.3V
V2 net3 GND DC 1.65V
**** begin user architecture code


.op
.control
set nobreak
set nomoremode
run
let power_val = v(vdd)*(-i(V1))
let current_val = (-i(V1))
echo 'POWER:' $&power_val
echo 'CURRENT:' $&current_val
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
