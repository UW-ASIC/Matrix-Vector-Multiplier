** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/TIAs/OpAmp_temp_opt/tb/OpAmp_TO_dc_gain_tb.sch
**.subckt OpAmp_TO_dc_gain_tb
**.ends
.end
