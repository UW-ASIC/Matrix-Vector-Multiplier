** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/TIAs/TIA_Balanced/tb/TIA_BAL_stability_analysis_tb.sch
**.subckt TIA_BAL_stability_analysis_tb
*  x1 -  TIA  IS MISSING !!!!
I0 net1 Iin DC 1u AC 1u
V1 net2 GND DC 3.3V
V2 net3 GND DC 1.65V
**** begin user architecture code


.ac dec 100 1 1G
.control
run
let gain_margin = 0
let phase_margin = 0
let unity_gain_freq = 0
let i = 0
while i < length(vdb(vout))
  if vdb(vout)[i] <= 0
    let unity_gain_freq = frequency[i]
    let phase_margin = 180 + vp(vout)[i]
    break
  end
  let i = i + 1
end
echo 'UNITY_GAIN_FREQ:' $&unity_gain_freq
echo 'PHASE_MARGIN:' $&phase_margin
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
