magic
tech sky130A
magscale 1 2
timestamp 1753657898
<< checkpaint >>
rect -541 1846 3457 3517
rect -541 1793 4276 1846
rect -541 1740 5617 1793
rect -1260 -1207 5617 1740
rect -1260 -1260 3457 -1207
rect -541 -1313 3457 -1260
<< error_p >>
rect 351 868 386 902
rect 352 849 386 868
rect 371 354 386 849
rect 405 815 440 849
rect 720 815 755 849
rect 405 354 439 815
rect 721 796 755 815
rect 1107 796 1160 797
rect 551 747 609 753
rect 551 713 563 747
rect 551 707 609 713
rect 551 437 609 443
rect 551 403 563 437
rect 551 397 609 403
rect 405 320 420 354
rect 740 301 755 796
rect 774 762 809 796
rect 1089 762 1160 796
rect 774 301 808 762
rect 1090 761 1160 762
rect 1107 727 1178 761
rect 1458 727 1493 761
rect 920 694 978 700
rect 920 660 932 694
rect 920 654 978 660
rect 920 384 978 390
rect 920 350 932 384
rect 920 344 978 350
rect 774 267 789 301
rect 1107 248 1177 727
rect 1459 708 1493 727
rect 1289 659 1347 665
rect 1289 625 1301 659
rect 1289 619 1347 625
rect 1289 331 1347 337
rect 1289 297 1301 331
rect 1289 291 1347 297
rect 1107 212 1160 248
rect 1478 195 1493 708
rect 1512 674 1547 708
rect 1512 195 1546 674
rect 1658 606 1716 612
rect 1658 572 1670 606
rect 1658 566 1716 572
rect 3199 553 3257 559
rect 3199 519 3211 553
rect 3199 513 3257 519
rect 4340 482 4398 488
rect 1658 278 1716 284
rect 1658 244 1670 278
rect 1658 238 1716 244
rect 1512 161 1527 195
rect 2810 118 2866 480
rect 4340 448 4352 482
rect 4340 442 4398 448
rect 2870 106 2926 420
rect 3199 225 3257 231
rect 3199 191 3211 225
rect 3199 185 3257 191
rect 4340 172 4398 178
rect 4340 138 4352 172
rect 4340 132 4398 138
use OpAmp  x1
timestamp 1753657898
transform 1 0 53 0 1 2371
box -53 -2371 4527 200
use sky130_fd_pr__cap_mim_m3_1_9C22PS  XC1
timestamp 0
transform 1 0 386 0 1 240
box -386 -240 386 240
use sky130_fd_pr__res_xhigh_po_5p73_J7EAP5  XR2
timestamp 0
transform 1 0 1458 0 1 1102
box -739 -1155 739 1155
<< end >>
