** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/Operational_Amplifiers/OpAmp_HighSpeed/tb/OpAmp_HS_dc_gain_tb.sch
**.subckt OpAmp_HS_dc_gain_tb
x1 vdd vout V- V+ net2 net1 OpAmp_HS
V1 net3 net4 DC 0.9V
V2 vdd GND DC 1.8V
V4 net2 net1 DC 0.7V
C1 vout GND 5p m=1
V3 V+ net3 DC 0V AC 1V
V5 V- net3 DC 0V
**** begin user architecture code


.ac dec 100 0.1 1G
.control
run
let dc_gain_val = vdb(vout)[0]
echo 'DC_GAIN:' $&dc_gain_val
let gbw_freq = 0
let i = 0
while i < length(vdb(vout))
  if vdb(vout)[i] <= 0
    let gbw_freq = frequency[i]
    break
  end
  let i = i + 1
end
echo 'GBW:' $&gbw_freq
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/omare/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  Operational_Amplifiers/OpAmp_HighSpeed/OpAmp_HS.sym # of pins=6
** sym_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/Operational_Amplifiers/OpAmp_HighSpeed/OpAmp_HS.sym
** sch_path: /home/omare/Documents/UWASIC/Matrix-Vector-Analog/analog/library/Operational_Amplifiers/OpAmp_HighSpeed/OpAmp_HS.sch
.subckt OpAmp_HS VDD Vout Vminus Vplus Vbias VSS
*.ipin Vplus
*.ipin Vminus
*.iopin VDD
*.iopin VSS
*.ipin Vbias
*.opin Vout
XM1 net2 Vminus net1 VSS sky130_fd_pr__nfet_01v8 L=0.18 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 Vplus net1 VSS sky130_fd_pr__nfet_01v8 L=0.18 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.18 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 Vbias VSS VSS sky130_fd_pr__nfet_01v8 L=0.18 W=100 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.40 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 Vout net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
XM7 Vout Vbias VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.GLOBAL VSS
.end
